module shiftLeft2bits(input logic[31:0] entrada, output logic [31:0] saida);

always_comb begin
	saida = entrada << 2;
end

endmodule: shiftLeft2bits